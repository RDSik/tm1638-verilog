// `define USE_HCW132_VARIANT_OF_TM1638_BOARD_CONTROLLER_MODULE
`define SPLIT_TM1638_DIO_INOUT_SIGNAL
// `define EMULATE_DYNAMIC_7SEG_ON_STATIC_WITHOUT_STICKY_FLOPS
`define NO_RESET_SYNCHRONIZER
